module rgmii_driver(
    input clk, rst,
    // RGMII signals
    inout [3:0] rgmii_txd,
    input rgmii_tx_ctl,
    input rgmii_rx_ctl,
    input [3:0] rgmii_rxd,
    output rgmii_rx_clk,
    output reg rst_n = 0,
    output reg [3:0] out = 0,
    output reg outclk = 0, 
    output reg done
);

`include "params.vh"

// RGMII Clock Skew
localparam RGMII_CLK_SKEW = 0; // Adjust this value as necessary

// RGMII clock is generated by the PHY
assign rgmii_rx_clk = clk; // Use system clock for simplicity

// RESET CONFIGURATION

// Similar to RMII, configure default settings after reset
localparam DEFAULT_MODE = 4'b0111; // Placeholder for default mode
localparam DEFAULT_PHYAD = 0;
localparam DEFAULT_NINTSEL = 1;

// Similar to RMII, set default values for RGMII signals after reset
assign rgmii_txd = rst_n ? 4'bz : DEFAULT_MODE;
assign rgmii_rx_ctl = rst_n ? 1'bz : DEFAULT_PHYAD;
assign rgmii_tx_ctl = rst_n ? 1'bz : DEFAULT_NINTSEL;

// RGMII does not require synchronization of signals

// RGMII PHY Interface State Machine
localparam STATE_IDLE = 0;
localparam STATE_WAITING = 1;
localparam STATE_PREAMBLE = 2;
localparam STATE_RECEIVING = 3;

reg [1:0] state = STATE_IDLE;

// Counter for RGMII clock skew
reg [3:0] rgmii_clk_count = 0;

always @(posedge clk) begin
    if (rst) begin
        rst_n <= 0;
        state <= STATE_IDLE;
        out <= 0;
        outclk <= 0;
        done <= 0;
        rgmii_clk_count <= 0;
    end else if (rst_n == 0 && rgmii_clk_count == RGMII_CLK_SKEW) begin
        rst_n <= 1;
    end else begin
        rgmii_clk_count <= rst_n ? 0 : (rgmii_clk_count + 1);
        case(state)
            STATE_IDLE:
                if (rgmii_rx_ctl)
                    state <= STATE_WAITING;
            STATE_WAITING:
                if (!rgmii_rx_ctl)
                    state <= STATE_IDLE;
                else if (rgmii_rxd == 4'b0001) // Preamble pattern detection
                    state <= STATE_PREAMBLE;
            STATE_PREAMBLE:
                if (!rgmii_rx_ctl)
                    state <= STATE_IDLE;
                else if (rgmii_rxd == 4'b1111) // End of preamble
                    state <= STATE_RECEIVING;
            STATE_RECEIVING:
                if (!rgmii_rx_ctl) begin
                    state <= STATE_IDLE;
                    outclk <= 0;
                    done <= 1; // Indicate frame reception completion
                end else begin
                    outclk <= 1;
                    out <= rgmii_rxd;
                end
        endcase
    end
end

endmodule
